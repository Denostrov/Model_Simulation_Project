radar format: 
x y z 
target format: 
x1 y1 z1 x2 y2 z2 x3 y3 z3  ...
max_load velocity
control center format:
x y z
launch silo format:
x y z
num_missile

Radars: 3
0 0 0
0 0 50
0 0 -50
Targets: 5
50 0 0 -50 0 0
5.0 5.0
50 0 25 -50 0 25
5.0 5.0
50 0 -25 -50 0 -25
5.0 5.0
50 0 50 -50 0 50
5.0 5.0
50 0 -50 -50 0 -50
5.0 5.0
ControlCenters: 1
-25 0 0
LaunchSilos: 2
-25 0 -50
4
-25 0 50
4

radar format: 
x y z 
target format: 
x1 y1 z1 x2 y2 z2 x3 y3 z3  ...
max_load velocity
control center format:
x y z
launch silo format:
x y z
num_missile

Radars: 5
60 0 -80
20 0 60
-60 0 40
-40 0 -50
0 0 -100
Targets: 8
100 20 -40 80 30 -60 60 20 -80
5 5
70 10 40 -50 20 10 40 20 70
5 4
60 20 100 30 20 0
5 4
40 40 -20 20 40 -80 -20 40 -80
5 4
-10 40 20 -40 20 30 -60 20 -10 -70 30 -30
5 4
-80 20 -10 -40 20 20 0 20 60
5 4
40 20 20 40 20 60
5 4
-60 10 -90 0 10 -40 -40 0 -40
5 4
ControlCenters: 1
0 0 -30
LaunchSilos: 3
80 0 0
6
-40 0 50
4
0 0 0
5
radar format: 
x y z 
target format: 
x1 y1 z1 x2 y2 z2 x3 y3 z3  ...
max_load velocity
control center format:
x y z
launch silo format:
x y z
num_missile

Radars: 2
0 0 -40
0 0 40
Targets: 20
50 10 -90 0 0 -40
5.0 5.0
50 10 -80 0 0 -40
5.0 3.0
50 10 -70 0 0 -40
5.0 5.0
50 10 -60 0 0 -40
5.0 3.0
50 10 -50 0 0 -40
5.0 5.0
50 10 -40 0 0 -40
5.0 3.0
50 10 -30 0 0 -40
5.0 5.0
50 10 -20 0 0 -40
5.0 3.0
50 10 -10 0 0 -40
5.0 5.0
50 10 0 0 0 -40
5.0 3.0
50 10 10 0 0 40
5.0 5.0
50 10 20 0 0 40
5.0 3.0
50 10 30 0 0 40
5.0 5.0
50 10 40 0 0 40
5.0 3.0
50 10 50 0 0 40
5.0 5.0
50 10 60 0 0 40
5.0 3.0
50 10 70 0 0 40
5.0 5.0
50 10 80 0 0 40
5.0 3.0
50 10 90 0 0 40
5.0 5.0
50 10 100 0 0 40
5.0 3.0
ControlCenters: 1
-25 0 0
LaunchSilos: 2
-25 0 -50
10
-25 0 50
10